--from SourceCode
library IEEE;
use IEEE.compoment;

entity test is port(..)
